* OPA172 - Rev. A
* Created by Ramon Jimenez, Paul Goedeke; August 01, 2018
* Created with Green-Williams-Lis Op Amp Macro-model Architecture
* Copyright 2018 by Texas Instruments Corporation
******************************************************
* MACRO-MODEL SIMULATED PARAMETERS:
******************************************************
* OPEN-LOOP GAIN AND PHASE VS. FREQUENCY  WITH RL, CL EFFECTS (Aol)
* UNITY GAIN BANDWIDTH (GBW)
* INPUT COMMON-MODE REJECTION RATIO VS. FREQUENCY (CMRR)
* POWER SUPPLY REJECTION RATIO VS. FREQUENCY (PSRR)
* DIFFERENTIAL INPUT IMPEDANCE (Zid)
* COMMON-MODE INPUT IMPEDANCE (Zic)
* OPEN-LOOP OUTPUT IMPEDANCE VS. FREQUENCY (Zo)
* OUTPUT CURRENT THROUGH THE SUPPLY (Iout)
* INPUT VOLTAGE NOISE DENSITY VS. FREQUENCY (en)
* INPUT CURRENT NOISE DENSITY VS. FREQUENCY (in)
* OUTPUT VOLTAGE SWING vs. OUTPUT CURRENT (Vo)
* SHORT-CIRCUIT OUTPUT CURRENT (Isc)
* QUIESCENT CURRENT (Iq)
* SETTLING TIME VS. CAPACITIVE LOAD (ts)
* SLEW RATE (SR)
* SMALL SIGNAL OVERSHOOT VS. CAPACITIVE LOAD
* LARGE SIGNAL RESPONSE
* OVERLOAD RECOVERY TIME (tor)
* INPUT BIAS CURRENT (Ib)
* INPUT OFFSET CURRENT (Ios)
* INPUT OFFSET VOLTAGE (Vos)
* INPUT COMMON-MODE VOLTAGE RANGE (Vcm)
* INPUT OFFSET VOLTAGE VS. INPUT COMMON-MODE VOLTAGE (Vos vs. Vcm)
* INPUT/OUTPUT ESD CELLS (ESDin, ESDout)
******************************************************
.subckt OPA172 IN+ IN- VCC VEE OUT
******************************************************
* MODEL DEFINITIONS:
.model BB_SW VSWITCH(Ron=50 Roff=1e12 Von=700e-3 Voff=0)
.model ESD_SW VSWITCH(Ron=50 Roff=1e12 Von=250e-3 Voff=0)
.model OL_SW VSWITCH(Ron=1e-3 Roff=1e9 Von=900e-3 Voff=800e-3)
.model OR_SW VSWITCH(Ron=10e-3 Roff=1e9 Von=1e-3 Voff=0)
.model R_NOISELESS RES(T_ABS=-273.15)
******************************************************


V_GRp       57 MID 60
V_GRn       58 MID -60
V_ISCp      51 MID 75
V_ISCn      52 MID -75
V_ORn       32 VCLP -1.75
V11         56 31 0
V_ORp       30 VCLP 1.75
V12         55 29 0
V4          45 OUT 0
VCM_MIN     79 VEE_B -100M
VCM_MAX     80 VCC_B -2
I_Q         VCC VEE 1.6M
I_OS        38 MID 6P
I_B         81 MID 8P
V_OS        87 21 164.1U
Xe_n        21 ESDp VNSE_0
C15         22 23 568.4P  
R55         23 22 R_NOISELESS 10K 
R56         MID 22 R_NOISELESS 9.342 
R54         MID 23 R_NOISELESS 1 
G_adjust2   23 MID 24 MID  -1
S11         ESDn ESDp ESDn ESDp  S_VSWITCH_1
S10         ESDp ESDn ESDp ESDn  S_VSWITCH_2
S5          VEE ESDp VEE ESDp  S_VSWITCH_3
S4          VEE ESDn VEE ESDn  S_VSWITCH_4
S2          ESDn VCC ESDn VCC  S_VSWITCH_5
S3          ESDp VCC ESDp VCC  S_VSWITCH_6
C28         25 MID 1P  
R75         26 25 R_NOISELESS 100 
C27         27 MID 1P  
R72         28 27 R_NOISELESS 100 
R74         MID 29 R_NOISELESS 1 
G11         29 MID 30 MID  -1
R73         31 MID R_NOISELESS 1 
G10         31 MID 32 MID  -1
R76         33 MID R_NOISELESS 1 
XVCCS_LIM_ZO 34 MID MID 33 VCCS_LIM_ZO_0
Xi_nn       ESDn MID FEMT_0
Xi_np       MID 21 FEMT_0
C25         35 MID 6.13F  
R69         MID 35 R_NOISELESS 1MEG 
G7          35 MID VSENSE MID  -1U
C20         CLAMP MID 50.1N  
R68         MID CLAMP R_NOISELESS 1MEG 
XVCCS_LIM_2 36 MID MID CLAMP VCCS_LIM_2_0
R44         MID 36 R_NOISELESS 1MEG 
XVCCS_LIM_1 37 38 MID 36 VCCS_LIM_1_0
R66         39 MID R_NOISELESS 1 
G6          39 MID 40 MID  -1
C23         41 MID 17.68P  
R65         40 41 R_NOISELESS 10K 
R64         40 42 R_NOISELESS 1.99MEG 
C26         39 34 636.6F  
R71         34 MID R_NOISELESS 2.5 
R70         34 39 R_NOISELESS 10K 
Rdc_1       42 MID R_NOISELESS 1 
G4          42 MID 43 MID  -590
C22         44 43 7.23U  
R51         43 MID R_NOISELESS 16.9 
R50         43 44 R_NOISELESS 10K 
Rdummy      MID 45 R_NOISELESS 1.65K 
Rx          45 33 R_NOISELESS 16.5K 
Rdc1        44 MID R_NOISELESS 1 
G_Aol_Zo    44 MID CL_CLAMP 45  -88
R62         MID 46 R_NOISELESS 106.7 
C21         46 47 4.974N  
R63         47 46 R_NOISELESS 100MEG 
G_adjust4   47 MID VEE_B MID  -937.5M
Rsrc3       MID 47 R_NOISELESS 1 
R57         MID 48 R_NOISELESS 148.1 
C16         48 49 159.2P  
R61         49 48 R_NOISELESS 100MEG 
G_adjust3   49 MID VCC_B MID  -675M
Rsrc2       MID 49 R_NOISELESS 1 
R48         MID 24 R_NOISELESS 93.42K 
C14         24 50 56.84F  
R49         50 24 R_NOISELESS 100MEG 
G_adjust1   50 MID ESDp MID  -1.071M
Rsrc1       MID 50 R_NOISELESS 1 
XIQp        VIMON MID MID VCC VCCS_LIMIT_IQ_0
XIQn        MID VIMON VEE MID VCCS_LIMIT_IQ_0
C_DIFF      ESDp ESDn 4P  
XCL_AMP     51 52 VIMON MID 53 54 CLAMP_AMP_LO_0
S8          CLAMP 55 CLAMP 55  S_VSWITCH_7
S9          56 CLAMP 56 CLAMP  S_VSWITCH_8
XGR_AMP     57 58 59 MID 60 61 CLAMP_AMP_HI_0
R39         57 MID R_NOISELESS 1T 
R37         58 MID R_NOISELESS 1T 
R42         VSENSE 59 R_NOISELESS 1M 
C19         59 MID 1F  
R38         60 MID R_NOISELESS 1 
R36         MID 61 R_NOISELESS 1 
R40         60 62 R_NOISELESS 1M 
R41         61 63 R_NOISELESS 1M 
C17         62 MID 1F  
C18         MID 63 1F  
XGR_SRC     62 63 CLAMP MID VCCS_LIM_GR_0
R35         53 MID R_NOISELESS 1 
R21         MID 54 R_NOISELESS 1 
R29         53 64 R_NOISELESS 1M 
R30         54 65 R_NOISELESS 1M 
C9          64 MID 1F  
C8          MID 65 1F  
XCL_SRC     64 65 CL_CLAMP MID VCCS_LIM_4_0
R22         51 MID R_NOISELESS 1T 
R20         MID 52 R_NOISELESS 1T 
XCLAWp      VIMON MID 66 VCC_B VCCS_LIM_CLAW+_0
XCLAWn      MID VIMON VEE_B 67 VCCS_LIM_CLAW-_0
R19         66 VCC_B R_NOISELESS 1K 
R16         66 68 R_NOISELESS 1M 
R13         VEE_B 67 R_NOISELESS 1K 
R17         69 67 R_NOISELESS 1M 
C6          69 MID 1F  
C5          MID 68 1F  
G2          VCC_CLP MID 68 MID  -1M
R15         VCC_CLP MID R_NOISELESS 1K 
G3          VEE_CLP MID 69 MID  -1M
R14         MID VEE_CLP R_NOISELESS 1K 
XCLAW_AMP   VCC_CLP VEE_CLP VOUT_S MID 70 71 CLAMP_AMP_LO_0
R26         VCC_CLP MID R_NOISELESS 1T 
R23         VEE_CLP MID R_NOISELESS 1T 
R25         70 MID R_NOISELESS 1 
R24         MID 71 R_NOISELESS 1 
R27         70 72 R_NOISELESS 1M 
R28         71 73 R_NOISELESS 1M 
C11         72 MID 1F  
C10         MID 73 1F  
XCLAW_SRC   72 73 CLAW_CLAMP MID VCCS_LIM_3_0
H2          28 MID V11 -1
H3          26 MID V12 1
C12         SW_OL MID 1P  
R32         74 SW_OL R_NOISELESS 100 
R31         74 MID R_NOISELESS 1 
XOL_SENSE   MID 74 27 25 OL_SENSE_0
S1          44 43 SW_OL MID  S_VSWITCH_9
H1          75 MID V4 1K
S7          VEE OUT VEE OUT  S_VSWITCH_10
S6          OUT VCC OUT VCC  S_VSWITCH_11
R12         MID 76 R_NOISELESS 1T 
R18         76 VOUT_S R_NOISELESS 100 
C7          VOUT_S MID 10P  
E5          76 MID OUT MID  1
C13         VIMON MID 1N  
R33         75 VIMON R_NOISELESS 100 
R11         MID 75 R_NOISELESS 1T 
R47         77 VCLP R_NOISELESS 100 
C24         VCLP MID 1P  
E4          77 MID CL_CLAMP MID  1
R46         MID CL_CLAMP R_NOISELESS 1K 
G9          CL_CLAMP MID CLAW_CLAMP MID  -1M
R45         MID CLAW_CLAMP R_NOISELESS 1K 
G8          CLAW_CLAMP MID 35 MID  -1M
R43         MID VSENSE R_NOISELESS 1K 
G15         VSENSE MID CLAMP MID  -1M
C4          37 MID 1F  
R10         37 78 R_NOISELESS 1M 
R9          MID 79 R_NOISELESS 1T 
R7          80 MID R_NOISELESS 1T 
R8          MID 78 R_NOISELESS 1 
XVCM_CLAMP  81 MID 78 MID 80 79 VCCS_EXT_LIM_0
E1          MID 0 82 0  1
R89         VEE_B 0 R_NOISELESS 1 
R6          83 VEE_B R_NOISELESS 1M 
C3          83 0 1F  
R60         82 83 R_NOISELESS 1MEG 
C1          82 0 1  
R5          82 0 R_NOISELESS 1T 
R59         84 82 R_NOISELESS 1MEG 
C2          84 0 1F  
R4          VCC_B 84 R_NOISELESS 1M 
R88         VCC_B 0 R_NOISELESS 1 
G17         VEE_B 0 VEE 0  -1
G16         VCC_B 0 VCC 0  -1
R67         85 81 R_NOISELESS 1K 
G1          81 85 48 46  -1M
R3          38 ESDn R_NOISELESS 1M 
R2          85 86 R_NOISELESS 1M 
R58         87 86 R_NOISELESS 1K 
G5          86 87 22 MID  -1
C_CMn       ESDn MID 4P  
C_CMp       MID ESDp 4P  
R53         ESDn MID R_NOISELESS 1T 
R52         MID ESDp R_NOISELESS 1T 
R1          IN- ESDn R_NOISELESS 250 
R34         IN+ ESDp R_NOISELESS 250 

.MODEL S_VSWITCH_1 VSWITCH (RON=50 ROFF=1T VON=700M VOFF=0)
.MODEL S_VSWITCH_2 VSWITCH (RON=50 ROFF=1T VON=700M VOFF=0)
.MODEL S_VSWITCH_3 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)
.MODEL S_VSWITCH_4 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)
.MODEL S_VSWITCH_5 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)
.MODEL S_VSWITCH_6 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)
.MODEL S_VSWITCH_7 VSWITCH (RON=10M ROFF=1T VON=1M VOFF=0)
.MODEL S_VSWITCH_8 VSWITCH (RON=10M ROFF=1T VON=1M VOFF=0)
.MODEL S_VSWITCH_9 VSWITCH (RON=1M ROFF=1T VON=900M VOFF=800M)
.MODEL S_VSWITCH_10 VSWITCH (RON=50 ROFF=1G VON=500M VOFF=100M)
.MODEL S_VSWITCH_11 VSWITCH (RON=50 ROFF=1G VON=500M VOFF=100M)

.ENDS OPA172
*
.SUBCKT VNSE_0  1 2
.PARAM FLW=1
.PARAM NLF=170
.PARAM NVR=6.2
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS VNSE_0 
*


.SUBCKT VCCS_LIM_ZO_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 4E3
.PARAM IPOS = 3.5E3
.PARAM INEG = -3.5E3
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT FEMT_0  1 2
.PARAM FLWF=1E-3
.PARAM NLFF=1.6
.PARAM NVRF=1.6
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
.ENDS FEMT_0 
*


.SUBCKT VCCS_LIM_2_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 3.68E-2
.PARAM IPOS = 0.50
.PARAM INEG = -0.50
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_1_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-4
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIMIT_IQ_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-3
G1 IOUT- IOUT+ VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
.ENDS
*


.SUBCKT CLAMP_AMP_LO_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=1
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT CLAMP_AMP_HI_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=10
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT VCCS_LIM_GR_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 1.2
.PARAM INEG = -1.2
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_4_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.26
.PARAM INEG = -0.26
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_CLAW+_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0, 1E-5)
+(23.65, 7.53E-4)
+(42.58, 1.14E-3)
+(60.97, 2.42E-3)
+(66.75, 2.87E-3)
+(76, 4.81E-3)
.ENDS
*


.SUBCKT VCCS_LIM_CLAW-_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0, 1E-5)
+(22.15, 1.2E-4)
+(40.77, 9.17E-4)
+(53.66, 1.56E-3)
+(67.77, 2.76E-3)
+(72.74, 3.46E-3)
+(76, 4.61E-3)
.ENDS
*


.SUBCKT VCCS_LIM_3_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.13
.PARAM INEG = -0.13
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT OL_SENSE_0  COM SW+ OLN  OLP
GSW+ COM SW+ VALUE = {IF((V(OLN,COM)>10E-3 | V(OLP,COM)>10E-3),1,0)}
.ENDS
*


.SUBCKT VCCS_EXT_LIM_0  VIN+ VIN- IOUT- IOUT+ VP+ VP-
.PARAM GAIN = 1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ENDS
*


